function Bool implies(Bool x, Bool y) = !x || y;
